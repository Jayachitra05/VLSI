class scoreboard;
  mailbox mail;
  transaction pkt;
  
  function new(mailbox mail);
    this.mail = mail;
  endfunction
  
  
