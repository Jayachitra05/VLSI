class adder_transaction;
  rand bit [3:0] a, b;  
  bit [3:0] y;         
endclass
