interface adder_if;
  logic [3:0] a, b;
  logic [3:0] y; 
endinterface
